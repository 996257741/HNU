module mux3_1(a,b,c,s,y);
    input [1:0] s;
	input [7:0] a,b,c;
	output reg[7:0] y;

always @(*) //alwaysģ���е��κ�һ�������źŻ��ƽ�����仯ʱ��������·���ģ�齫��ִ��
    begin
    if(s==2'b00) y=a;
    else if(s==2'b01) y=b;
    else if(s==2'b10) y=c;
    else y=a;
    end
endmodule